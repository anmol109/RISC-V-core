module riscv_alu
(
    // Inputs
input clk,rst,
input is_beq,is_bne,is_blt,is_bge,is_bltu,is_bgeu,
is_add,
is_addi,
is_slti,
is_or,
is_ori,
is_xor,
is_xori,
is_and,
is_andi,
is_sub,
is_sltiu,
is_slli,
is_srli,
is_srai,
is_sll,
is_slt,
is_sltu,
is_srl,
is_sra,
is_lui,
is_auipc,
is_jal,
is_jalr,
is_jump,
is_lb,
is_lh,
is_lw,
is_lbu,
is_lhu,
is_sb,
is_sh,
is_sw,
is_ecall,
    input  [ 31:0]  alu_a
    ,input  [ 31:0]  alu_b

    // Outputs
    ,output [ 31:0]  alu_p_o
);
reg[31:0] result,a_r,b_r;

always@(posedge clk) begin
if(is_add || is_addi) //add instruction
result=alu_a+alu_b;
else if(is_sub)// sub instr
result=alu_a-alu_b;
else if(is_or || is_ori) // or instr
result=alu_a||alu_b;
else if(is_xor||is_xori) //xor instr
result=alu_a^alu_b;
else if(is_and||is_andi) //and instr
result=alu_a&alu_b;
else if(is_sll||is_slli) //logical left shift
result=alu_a<<alu_b;
else if(is_srl||is_srli)
result=alu_a>>alu_b; //logical right shift
else if(is_sra||is_srai)
result=alu_a>>>alu_b; //arithmetic right shift
else if(is_sltiu||is_sltu)begin
	if(alu_a>alu_b)
		result=alu_b;
	else 
		result=alu_a;
end
else if(is_slt||is_slti) begin
	if((alu_a==1'b1)&&(alu_b==1'b1))begin
		if(alu_a<alu_b)
			result=alu_b;
		else
			result=alu_a;
	end
	else begin
		a_r[30:0]=alu_a[30:0];
		b_r[30:0]=alu_b[30:0];
		a_r[31]=~alu_a[31];
		b_r[31]=~alu_b[31];
		if(a_r<b_r)
			result=alu_a;
		else
			result=alu_b;
	end
end
else
result=32'dx;
end




assign alu_p_o = result;

endmodule
