module rv_top();


